* fogor

* R30 V15_P V15_PF 0.00001
* R31 V15_N V15_NF 0.00001

.SUBCKT FERRITE_22U 1 3
R1 1 2 0.35
L1 2 3 22u
C1 1 3 1.3p
.ENDS

.SUBCKT LQM21FN4R7N00L 1 3
R1 1 2 0.3
L1 2 3 4.7u
C1 1 3 1.3p
.ENDS

.SUBCKT POWER
X1 V15_P 0 C0603C104K5RAC
X2 0 V15_N C0603C104K5RAC
X3 V15_P 0 C_100U
X4 0 V15_N C_100U

X5 V15_P V15_PF LQM21FN4R7N00L
X6 V15_N V15_NF LQM21FN4R7N00L

X10 V15_PF 0 C_100U
X11 0 V15_NF C_100U
X12 V15_PF 0 C_100U
X13 0 V15_NF C_100U
X14 V15_PF 0 C_100U
X15 0 V15_NF C_100U

X16 V15_PF 0 C0603C104K5RAC
X17 0 V15_NF C0603C104K5RAC

* R10 V15_PF 0 1000
* R11 V15_NF 0 1000

* v4000 V33 0 dc 3.3

* V334 V33 0 dc 3.3

X3 V15_PF 0 V33 REG33
R1 V33 V_CPU 0.001

* C931 V33 0 10m
*C932 V15_PF 0 10m
X100 V33 0 C_100U
*X101 V33 0 C_100U
* C100 V33 0 2.5p
* X101 V33A 0 C_100U
* X101 V33 0 C_100U
X110 V33 0 C0603C104K5RAC
X111 V33 0 C1206C104K2RAC
X112 V33 0 C1206C104K2RAC
* X113 V33A 0 C1206C104K2RAC

X120 V_CPU 0 C0603C104K5RAC
X121 V_CPU 0 C0603C104K5RAC

R2 V15_PF V15_NF 100k

* v1 V33 0 dc 3.3
* v2 VOFFSET 0 dc 1.65

R30 V33 VOFFSET 1k
R31 VOFFSET 0 1k
X300 VOFFSET 0 C0603C104K5RAC
* C300 VOFFSET 0 10m

R50 V33 V33A 0.001
* T1 V33 0 V33A 0 Z0=51 TD=0.56n

* X200 V33 V33A FERRITE_22U
* R200 V33 V33A 0.001
X201 V33A 0 C0603C104K5RAC
*X202 V33A 0 C_100U
* X202 V33A 0 C0603C104K5RAC
* X203 V33A 0 C0603C104K5RAC
*X204 V33A1 0 C0603C104K5RAC
* X202 V33A 0 C0603C104K5RAC

R202 V33A 0 825
.ENDS

.SUBCKT MFC 1 2 3 5
G1 3 4 1 2 3.5e-3
C1 3 4 84.04n
R1 3 4 10G
G2 2 1 3 4 3.5e-3
R2 4 5 0.01
.ENDS

.SUBCKT VEL_IN VIN VOUT V33 VOFFSET VP VN XGND
* measurement resistor
R1 VIN XGND 47

* RFI filter
R2 VIN V1 1k
C1 V1 XGND 1n

* Stage 1: +20 dB
R3 XGND V2F 10k
R4 V2F V2 100k
X1 V1 V2F VP VN V2 TL074NEW

R100 V2 V3 0.01

* Stage 2: +20 dB
R5 V3 V3F 10k
R6 V3F V4 100k
X3 1 V3F VP VN V4 TL074NEW
* X3 1 V3F VP VN V4 LM224

R8 VOFFSET 1 100k
R9 1 XGND 10k

* ADC: filter
*R7 V4 VOUT 1k
*C3 VOUT XGND 1n

R7 V4 VOUT 47
C3 VOUT XGND 1n
*C3 VOUT XGND 100n

* v1 VZZ XGND dc 3
* X10 XGND VOUT VP VN VOUT TL074NEW
* R101 VOUT XGND 10k
.ENDS

.SUBCKT A_IN VIN VOUT V33 VOFFSET VP VN XGND
* RFI filter
R1 VIN V1 1k
C1 V1 XGND 1n

R2 V1 V2 1000k
R3 V2 XGND 100k

X1 V2 V3 VP VN V3 TL074NEW

R4 V3 V4F 100k
R5 V4F V4 10k
X2 1 V4F VP VN V4 TL074NEW

R6 VOFFSET 1 10k
R7 1 XGND 100k

* ADC: filter
* R6 VOUT 0 1k
R9 V4 VOUT 1k
C3 VOUT XGND 1n
.ENDS

*
* PWM-based DAC
* Input: 3.3V peak-to-peak, +4.35 dB peak
* Output: line out, -10 dB nominal
* Bandwidth: 
*
.SUBCKT DAC VIN VOUT V33 XGND
R1 VIN V1 1k
X1 V1 XGND C0603C104K5RAC

R2 V1 V2 1k
* C2 V2 XGND 100n
X2 V2 XGND C0603C104K5RAC
* X2 V2 XGND C0603C104K5RAC
* C1 V2 XGND 10n

R3 V2 V33 1k
R4 V2 XGND 1k

* C1 V2 VOUT 100u
* X3 V2 VOUT C0603C104K5RAC
C3 V2 VOUT 100u
*R10 V2 VOUT 1
R5 VOUT XGND 1meg

* R6 VOUT XGND 47
.ENDS

.SUBCKT DAC4 VIN VOUT V33 XGND
R1 VIN V1 1k
* X1 V1 XGND C0603C104K5RAC
R2 V1 V2 1k

R33 V1 0 10meg

*R3 V2 V33 1k
* R4 V2 XGND 1k

C3 V2 VOUT 100u
R5 VOUT XGND 1k
X2 VOUT XGND C0603C104K5RAC
.ENDS


.SUBCKT DAC3 VIN VOUT V33 XGND
R1 VIN V1 220
X1 V1 XGND C0603C104K5RAC
R2 V1 V2 220

R33 V1 0 10meg

*R3 V2 V33 1k
*R4 V2 XGND 1k

C3 V2 VOUT 10u
R5 VOUT XGND 100
X2 VOUT XGND C0603C104K5RAC
.ENDS

.SUBCKT LINEIN VIN VOUT V33 XGND
R1 VIN V1 10k
*C1 V1 XGND 1n

R2 VIN V2 10k
* R30 V2 VOUT 0.001
X2 V2 VOUT C0603C104K5RAC

R3 VOUT V33 100k
R30 VOUT V33 100k
* R31 VOUT V33 100k
R4 VOUT XGND 100k

* C2 VOUT XGND 1n
X3 VOUT XGND C0603C104K5RAC
.ENDS

.SUBCKT LINEINX VIN VOUT V33 XGND
R1 VIN V1 10k
*C1 V1 XGND 1n

R2 VIN V2 10k
* R30 V2 VOUT 0.001
X2 V2 VOUT C0603C104K5RAC

R3 VOUT V33 1000k
R4 VOUT XGND 1000k

C2 VOUT XGND 1n
.ENDS

.SUBCKT TRAFO p1 p2 s1 s2 N=1 L=1
L1 p1 p2 {L}
L2 s1 s2 {N*N*L}
K1 L1 L2 1
.ENDS

.SUBCKT RECOVERY MFC V_PLUS V_MINUS XGND
C100 MFC XGND 110u
L100 MFC XGND 10.235m
* L100 MFCX XGND 3.26

* X1 MFCX XGND MFC XGND TRAFO N=10 L=3.26

* D10 XGND MFC LL4148

D1 MFC V_PLUS LL4148
C1 V_PLUS XGND 100u
D2 XGND V_PLUS LL4148
D3 V_PLUS V1 LL4148
D4 V1 V2 LL4148
D5 V2 V3 LL4148
D6 V3 V4 LL4148
D7 V4 XGND LL4148

*v1 V_PLUS XGND dc 3.3
*v2 V_MINUS XGND dc 0

D11 V_MINUS MFC LL4148
C11 V_MINUS XGND 100u
D12 V_MINUS XGND LL4148
D13 XGND V1 LL4148
D14 V1 V2 LL4148
D15 V2 V3 LL4148
D16 V3 V4 LL4148
D17 V4 V_MINUS LL4148
.ENDS

.SUBCKT OUTSW MFC POS NEG V_PLUS V_MINUS V33 V15 VN15 XGND
R30 POS Q1B 10k
R32 Q1B XGND 10k
Q1 Q1C Q1B XGND BC847

R27 Q1C Q2B 10k
R28 Q2B V15 10k
Q2 Q2C Q2B V15 BC857

R23 Q2C Q3G 47
* FIXME
R24 Q2C 0 2.2k
X3 Q3D Q3G V_MINUS FQD12N20L
D4 MFC Q3D LL4148

* v1 V_MINUS 0 dc -3.3
* v2 V_PLUS 0 dc 3.3

*v1 V_MINUS 0 dc 0
*v2 V_PLUS 0 dc 0

R34 NEG Q4B 10k
R36 Q4B V33 10k
Q4 Q4C Q4B V33 BC857

R39 Q4C Q6B 10k
R40 Q6B VN15 10k
Q6 Q6C Q6B VN15 BC847

R26 Q6C Q5G 47
* FIXME
R25 Q6C 0 2.2k
X5 Q5D Q5G V_PLUS FQD7P20
D5 Q5D MFC LL4148
.ENDS
