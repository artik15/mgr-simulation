*foo

* TL074 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 06/16/89 AT 13:08
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TL074    1 2 3 4 55
*
  C1   11 12 3.498E-12
  C2    6  7 15.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 4.715E6 -5E6 5E6 5E6 -5E6
  GA    6  0 11 12 282.8E-6
  GCM   0  6 10 99 8.942E-9
  ISS   3 10 DC 195.0E-6
  HLIM 90  0 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100.0E3
  RD1   4 11 3.536E3
  RD2   4 12 3.536E3
  RO1   8  5 150
  RO2   7 99 150
  RP    3  4 2.143E3
  RSS  10 99 1.026E6
  VB    9  0 DC 0
  VC    3 53 DC 2.200
  VE   54  4 DC 2.200
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=15.00E-12 BETA=270.1E-6 VTO=-1)
  
  ROUT   5 55 0.0001
.ENDS

.SUBCKT TL074NEW    1 2 3 4 55
*
  C1   11 12 3.498E-12
  C2    6  7 15.00E-12
*   C2    6  7 15.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99 1000 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 4.715E6 -5E6 5E6 5E6 -5E6
  GA    6 1000 11 12 282.8E-6
  GCM   1000  6 10 99 8.942E-9
  ISS   3 10 DC 195.0E-6
  HLIM 90  1000 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6 9 100.0E3
  RD1   4 11 3.536E3
  RD2   4 12 3.536E3
  RO1   8  5 150
  RO2   7 99 150
  RP1    3  1000 1.0715E3
  RP2    1000  4 1.0715E3
  RSS  10 99 1.026E6
  VB    9 1000 DC 0
  VC    3 53 DC 2.200
  VE   54  4 DC 2.200
  VLIM  7  8 DC 0
  VLP  91  1000 DC 25
  VLN   1000 92 DC 25
.MODEL DX D(IS=800.0E-18 KF=1.5e-11)
* .MODEL DX D(IS=800.0E-18 KF=1.5e-11)
.MODEL JX PJF(IS=15.00E-12 BETA=270.1E-6 VTO=-1)

  RXX 0 1000 0.001
  
  ROUT   5 55 0.0001
.ENDS

.SUBCKT REG33 IN ADJ OUT
v1 1 IN dc 8
x1 1 ADJX OUT LM317
v2 ADJ ADJX dc -2.05
.ENDS

.SUBCKT LM317 in adj out
* PEI 08/98 p62
J1 in out 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL .2
Q4 8 5 7 QPL .1
Q5 81 8 out QNL .2
Q6 out 81 10 QPL .2
Q7 12 81 13 QNL .2
*Q8 10 5 11 QPL .2
Q8 10A 5 11 QPL .2
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL .2
Q11 16 14 15 QNL .2 OFF
Q12 out 20 16 QPL .2
Q13 in 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 out 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 out 24 QNL .2
Q18 22 22 16 QPL .2
Q19 22 out 241 QNL .2
Q20 out 25 16 QPL .2
Q21 25 26 out QNL .2
Q22A 35 35 in QPL .2
Q22B 16 35 in QPL .2
Q23 35 16 30 QNL .2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 in 31 41 QNL 5
Q26 in 41 32 QNL 50
D1 out 4 DZ
D2 33 in DZ
D3 29 34 DZ
R1 in 6 310
R2 in 7 310
R3 in 11 190
R4 in 17 82
R5 in 18 5.6K
R6 4 8 100K
R7 8 81 130
*R8 10 12 12.4K
R8 10A 12 12.4K
R9 9 out 180
R10 13 out 4.1K
R11 14 out 5.8K
R12 15 out 72
R13 20 out 5.1K
R14 adj 24 12K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 130
R19 16 31 370
R20 26 27 13K
R21 27 40 400
R22 out 41 160
R23 33 34 18K
R24 28 29 160
R25 28 32 3
R26 32 out .1
C1 21 out 30PF
C2 21 adj 30PF
C3 25 26 5PF
CBS1 5 out 2PF
CBS2 35 out 1PF
CBS3 22 out 1PF
.MODEL JN NJF (BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN (EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS
+ CJE=2PF CJC=1PF VAF=100 IS=1E-22 NF=1.2)
.MODEL QPL PNP (BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50
+ IS=1E-22 NF=1.2)
.ENDS LM317

.SUBCKT L1U5 1 3
L1 1 2 1.5u
R1 2 3 0.45
C1 1 3 20p
.ENDS

.SUBCKT C0603C104K5RAC 1 6
* Temp@ 25�C, Bias@ 0Vdc , Center Freq@ 1.000MHz
* KEMET Model RLC Cerm.JPG / Spice Version 3.9.5 
L1  1 2 99.50E-12
L2  2 3 1.89E-09
R1  3 4 139.41E-03
C1  4 6 91.00E-09
R2  2 5 10.6
C2  5 6 4.10E-12
R3  1 6 10.000E+09
.ENDS

.SUBCKT C_100U 1 4
L1  1 2 10n
R1  2 3 0.5
C1  3 4 100e-6
R2  1 4 1000k
.ENDS

.SUBCKT LM224    1   2  99  50  28
*
*Features:
*Eliminates need for dual supplies
*Large DC voltage gain =             100dB
*High bandwidth =                     1MHz
*Low input offset voltage =            2mV
*Wide supply range =        +-1.5V to +-16V
*
*NOTE: Model is for single device only and simulated
*      supply current is 1/4 of total device current.
*      Output crossover distortion with dual supplies
*      is not modeled.
*
****************INPUT STAGE**************
*
IOS 2 1 3N
*^Input offset current
R1 1 3 500K
R2 3 2 500K
I1 99 4 100U
R3 5 50 517
R4 6 50 517
Q1 5 2 4 QX
Q2 6 7 4 QX
*Fp2=1.2 MHz
C4 5 6 128.27P
*
***********COMMON MODE EFFECT***********
*
I2 99 50 75U
*^Quiescent supply current
EOS 7 1 POLY(1) 16 49 2E-3 1
*Input offset voltage.^
R8 99 49 60K
R9 49 50 60K
*
*********OUTPUT VOLTAGE LIMITING********
V2 99 8 1.63
D1 9 8 DX
D2 10 9 DX
V3 10 50 .635
*
**************SECOND STAGE**************
*
EH 99 98 99 49 1
G1 98 9 POLY(1) 5 6 0 9.8772E-4 0 .3459
*Fp1=7.86 Hz
R5 98 9 101.2433MEG
C3 98 9 200P
*
***************POLE STAGE***************
*
*Fp=2 MHz
G3 98 15 9 49 1E-6
R12 98 15 1MEG
C5 98 15 7.9577E-14
*
*********COMMON-MODE ZERO STAGE*********
*
*Fpcm=10 KHz
G4 98 16 3 49 5.6234E-8               
L2 98 17 15.9M
R13 17 16 1K
*
**************OUTPUT STAGE**************
*
F6 50 99 POLY(1) V6 300U 1
E1 99 23 99 15 1
R16 24 23 17.5
D5 26 24 DX
V6 26 22 .63V
R17 23 25 17.5
D6 25 27 DX
V7 22 27 .63V
V5 22 21 0.27V
D4 21 15 DX
V4 20 22 0.27V
D3 15 20 DX
L3 22 28 500P
RL3 22 28 100K
*
***************MODELS USED**************
*
.MODEL DX D(IS=1E-15)
.MODEL QX PNP(BF=1.111E3)
.ENDS


** Standard Linear Ics Macromodels, 1993. 
** CONNECTIONS :
* 1 INVERTING INPUT
* 2 NON-INVERTING INPUT
* 3 OUTPUT
* 4 POSITIVE POWER SUPPLY
* 5 NEGATIVE POWER SUPPLY
.SUBCKT TL07x 2 1 4 5 3
**********************************************************
.MODEL MDTH D IS=1E-8 KF=5.306587E-14 CJO=10F
* INPUT STAGE
CIP 2 5 1.000000E-12
CIN 1 5 1.000000E-12
EIP 10 5 2 5 1
EIN 16 5 1 5 1
RIP 10 11 1.130435E+00
RIN 15 16 1.130435E+00
RIS 11 15 2.476554E-01
DIP 11 12 MDTH 400E-12
DIN 15 14 MDTH 400E-12
VOFP 12 13 DC 0
VOFN 13 14 DC 0
IPOL 13 5 2.300000E-04
CPS 11 15 4.091333E-08
DINN 17 13 MDTH 400E-12
VIN 17 5 3.000000e+00
DINR 15 18 MDTH 400E-12
VIP 4 18 0.000000E+00
FCP 4 5 VOFP 6.096957E+00
FCN 5 4 VOFN 6.096957E+00
* AMPLIFYING STAGE
FIP 5 19 VOFP 8.217391E+02
FIN 5 19 VOFN 8.217391E+02
RG1 19 5 1.112645E+06
RG2 19 4 1.112645E+06
CC 19 29 1.300000E-08
HZTP 30 29 VOFP 7.743183E+02
HZTN  5 30 VOFN 7.743183E+02
DOPM 19 22 MDTH 400E-12
DONM 21 19 MDTH 400E-12
HOPM 22 28 VOUT 3.750000E+03
VIPM 28 4 1.500000E+02
HONM 21 27 VOUT 3.750000E+03
VINM 5 27 1.500000E+02
EOUT 26 23 19 5 1
VOUT 23 5 0
ROUT 26 3 9.384786E+01
COUT 3 5 1.000000E-12
DOP 19 25 MDTH 400E-12
VOP 4 25 3.259753E+00
DON 24 19 MDTH 400E-12
VON 24 5 3.259753E+00
.ENDS; TL07x

.SUBCKT C1206C104K2RAC 1 6
* Temp@ 25�C, Bias@ 0Vdc , Center Freq@ 1.000MHz
* KEMET Model RLC Cerm.JPG / Spice Version 3.9.5 
L1  1 2 99.50E-12
L2  2 3 1.89E-09
R1  3 4 67.98E-03
C1  4 6 91.00E-09
R2  2 5 5.6
C2  5 6 4.20E-12
R3  1 6 10.000E+09
.ENDS

*$
**************** Power Discrete MOSFET Electrical Circuit Model *****************
** Product Name: FQD12N20LTM
** 200V, 9.0A, 280mohm N-Channel QFET
** Model Type: BSIM3V3
**-------------------------------------------------------------------------------
.SUBCKT FQD12N20L 2 1 3    
*Nom Temp=25 deg C
Dbody 7 5    DbodyMOD
Dbreak 5 11  DbreakMOD
Ebreak 11 7 17 7 220
Lgate 1 9    1.183e-9
Ldrain 2 5   1.440e-9
Lsource 3 7  9.664e-10
RLgate 1 9   11.83
RLdrain 2 5  14.4
RLsource 3 7 9.66
Rgate 9 6    0.5
It 7 17      1
Rbreak 17 7  RbreakMOD 1
.MODEL RbreakMOD RES (TC1=9.18e-4 TC2=-1.13e-6)
.MODEL DbodyMOD D (IS=1.15e-12  N=1.0    RS=1.82e-2  TRS1=1.85e-3  TRS2=1.82e-7 
+ CJO=7.84e-10     M=0.66       VJ=0.46  TT=1.35e-7  XTI=3         EG=1.14)
.MODEL DbreakMOD D (RS=100e-3 TRS1=1.0e-3 TRS2=1e-6)
Rdrain 5 16 RdrainMOD 0.19
.MODEL RdrainMOD RES (TC1=7.62e-3 TC2=1.75e-5)
M_BSIM3 16 6 7 7 Bsim3 W=1.23 L=2.0e-6 NRS=1
.MODEL Bsim3 NMOS (LEVEL=49 VERSION=3.1 MOBMOD=3 CAPMOD=2 PARAMCHK=1 NQSMOD=0
+ TOX=500e-10     XJ=1.4e-6      NCH=1.23e17      
+ U0=700          VSAT=1.0e5     DROUT=1.0     
+ DELTA=0.1       PSCBE2=0       RSH=2.59e-2    
+ VTH0=1.75       VOFF=-0.1      NFACTOR=1.1
+ LINT=4.25e-7    DLC=4.25e-7    FC=0.5
+ CGSO=1.00e-15   CGSL=0         CGDO=2.05e-15 
+ CGDL=1.18e-9    CJ=0           CF=0
+ CKAPPA=0.2      KT1=-1.45      KT2=0
+ UA1=8.8e-9      NJ=10)
.ENDS
*$
********************* Power Discrete MOSFET Thermal Model **********************
** Package: D-PAK
**------------------------------------------------------------------------------
.SUBCKT FQD12N20L_Thermal TH TL
CTHERM1 TH 6 2.41e-4
CTHERM2 6 5  4.80e-3
CTHERM3 5 4  9.80e-3
CTHERM4 4 3  1.30e-2
CTHERM5 3 2  4.00e-2
CTHERM6 2 TL 1.20e-1 
RTHERM1 TH 6 1.96e-2
RTHERM2 6 5  6.76e-2
RTHERM3 5 4  7.98e-2
RTHERM4 4 3  1.83e-1
RTHERM5 3 2  5.99e-1
RTHERM6 2 TL 1.33e+0
.ENDS FQD12N20L_Thermal 
**------------------------------------------------------------------------------
** Creation: Jun.-15-2017   Rev.: 2.0
** ON Semiconductor
*$

.MODEL BC847 NPN
+     IS = 1.822E-14 
+     NF = 0.9932 
+     ISE = 2.894E-16 
+     NE = 1.4 
+     BF = 324.4 
+     IKF = 0.109 
+     VAF = 82 
+     NR = 0.9931 
+     ISC = 9.982E-12 
+     NC = 1.763 
+     BR = 8.29 
+     IKR = 0.09 
+     VAR = 17.9 
+     RB = 10 
+     IRB = 5E-06 
+     RBM = 5 
+     RE = 0.649 
+     RC = 0.7014 
+     XTB = 0 
+     EG = 1.11 
+     XTI = 3 
+     CJE = 1.244E-11 
+     VJE = 0.7579 
+     MJE = 0.3656 
+     TF = 4.908E-10 
+     XTF = 9.51 
+     VTF = 2.927 
+     ITF = 0.3131 
+     PTF = 0 
+     CJC = 3.347E-12 
+     VJC = 0.5463 
+     MJC = 0.391 
+     XCJC = 0.6193 
+     TR = 9E-08 
+     CJS = 0 
+     VJS = 0.75 
+     MJS = 0.333 
+     FC = 0.979

.MODEL BC857 PNP
+     IS = 2.014E-14 
+     NF = 0.9974 
+     ISE = 6.578E-15 
+     NE = 1.45 
+     BF = 315.3 
+     IKF = 0.079 
+     VAF = 39.15 
+     NR = 0.9952 
+     ISC = 1.633E-14 
+     NC = 1.15 
+     BR = 8.68 
+     IKR = 0.09 
+     VAR = 9.5 
+     RB = 10 
+     IRB = 5E-06 
+     RBM = 5E-06 
+     RE = 0.663 
+     RC = 0.718 
+     XTB = 0 
+     EG = 1.11 
+     XTI = 3 
+     CJE = 1.135E-11 
+     VJE = 0.7071 
+     MJE = 0.3808 
+     TF = 6.546E-10 
+     XTF = 5.387 
+     VTF = 6.245 
+     ITF = 0.2108 
+     PTF = 0 
+     CJC = 6.395E-12 
+     VJC = 0.4951 
+     MJC = 0.44 
+     XCJC = 0.6288 
+     TR = 5.5E-08 
+     CJS = 0 
+     VJS = 0.75 
+     MJS = 0.333  
+     FC = 0.9059
*

********* Discrete Diode Electrical Parameters *********
** Package: OSD80
** LL4148 Small Signal Diode
**------------------------------------------------------
.MODEL LL4148 D
+ IS=3.6e-9       RS=0.03622    N=2.0   
+ ISR=7.208e-9    NR=2.0        CJO=8.68e-13
+ M=0.021         VJ=0.6506     FC=0.5
+ TT=3.812e-9     BV=100.5      IBV=1.0e-4
+ EG=1.02         XTI=3
**------------------------------------------------------
** Creation: Jan.-03-2012   Rev: 0.0
** Fairchild Semiconductor

*FQD7P20 200V P-CHANNEL DMOSFET ELECTRICAL PARAMETERS
*------------------------------------------------------------------------------------
.SUBCKT  FQD7P20   20  10  30
.param TEMP = 27
Rg     10    1    1
M1      2    1    3    3    DMOS    L=1u   W=1u
.MODEL DMOS PMOS (VTO={-3.9*(-0.00088*TEMP+1.022)} KP={4.4*(-0.00012*TEMP+1.003)} 
+ THETA=0.04    VMAX=1.52E5   LEVEL=3)
Cgs 1   3   680P
Rd  20  4   236m   TC=0.00083
Dds 4   3   DDS
.MODEL DDS D(BV={200*(0.0008*TEMP+0.98)}  M=0.5      CJO=115p   VJ=0.8)
Dbody   20  3   DBODY
.MODEL DBODY D(IS=1.2E-13    N=1.05     RS=96.3m    EG=1.17    TT=180n)
Ra 4    2   110m   TC=0.00083
Rs 3    5   11m    
Ls 5    30  1.0n
M2 1    8   6    6   INTER
E2 8    6   4    1   2
.MODEL INTER PMOS (VTO=0   KP=10   LEVEL=1)
Cgdmax  7  4    925P
Rcgd    7  4    10meg
Dgd     4  6    DGD
Rdgd    4  6    10meg
.MODEL DGD D(M=0.74   CJO=925P    VJ=0.62)
M3      7  9  1  1  INTER
E3      9  1  4  1  -2
.ENDS FQD7P20
*-------------------------------------------------------------------------------------
*FAIRCHILD      CASE: D-PAK      PID: FQD7P20 
*NOV-18-2000 CREATION  
*.SUBCKT COIL 1 3
*L1 1 2 2.2m
*R1 2 3 1.6
*C1 1 3 61p
*.ENDS

.SUBCKT COILX 1 3
L1 1 2 1m
R1 2 3 3.85
C1 1 3 20p
.ENDS

.SUBCKT RC5256 1 3
L1 1 2 500u
R1 2 3 0.26
C1 1 3 52p
.ENDS

.SUBCKT RC5258 1 3
L1 1 2 1000u
R1 2 3 0.55
C1 1 3 60p
.ENDS

.SUBCKT COIL2 1 6
X1 1 2 RC5256
X2 2 3 RC5256
X3 3 4 RC5256
X4 4 5 RC5256
X5 5 6 RC5256
.ENDS

.SUBCKT COILXX 1 5
X1 1 2 RC5258
X2 2 3 RC5258
X3 3 4 RC5258
X4 4 5 RC5258
.ENDS

.SUBCKT COIL5 1 3
L1 1 2 30m
R1 2 3 2.7
C1 1 3 33p
.ENDS

.SUBCKT COILOLD 1 3
L1 1 2 2.5e-2
R1 2 3 7.5e-1
C1 1 3 2.3e-11
.ENDS
